module interleaver ();


endmodule